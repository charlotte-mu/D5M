module TOP(

);


endmodule
