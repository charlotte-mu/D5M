module D5M_rom(
	input [7:0] address,
	output [15:0] data_out
);
reg [15:0]rom[255:0];
assign data_out = rom[address];
initial
begin
		rom[0]   	<= 16'h1801;
		rom[1]   	<= 16'h0036;
		rom[2]   	<= 16'h0010;
		rom[3]   	<= 16'd1079;
		rom[4]   	<= 16'd1919;
		rom[5]   	<= 16'h0;
		rom[6]   	<= 16'h0019;
		rom[7]   	<= 16'h1f82;
		rom[8]   	<= 16'h0;
		rom[9]   	<= 16'h0797;
		rom[10]   	<= 16'h0;
		rom[11]   	<= 16'h0;
		rom[12]   	<= 16'h0;
		rom[13]   	<= 16'h0;
		rom[14]   	<= 16'h0;
		rom[15]   	<= 16'h0;
		rom[16]   	<= 16'h0050;
		rom[17]   	<= 16'h6404;
		rom[18]   	<= 16'h0;
		rom[19]   	<= 16'h0;
		rom[20]   	<= 16'h0036;
		rom[21]   	<= 16'h0010;
		rom[22]   	<= 16'h0;
		rom[23]   	<= 16'h0;
		rom[24]   	<= 16'h0;
		rom[25]   	<= 16'h0;
		rom[26]   	<= 16'h0;
		rom[27]   	<= 16'h0;
		rom[28]   	<= 16'h0;
		rom[29]   	<= 16'h0;
		rom[30]   	<= 16'h4006;
		rom[31]   	<= 16'h0;
		rom[32]   	<= 16'h0040;
		rom[33]   	<= 16'h0;
		rom[34]   	<= 16'h0;
		rom[35]   	<= 16'h0;
		rom[36]   	<= 16'h0002;
		rom[37]   	<= 16'h0;
		rom[38]   	<= 16'h0;
		rom[39]   	<= 16'h000b;
		rom[40]   	<= 16'h0;
		rom[41]   	<= 16'h0481;
		rom[42]   	<= 16'h1086;
		rom[43]   	<= 16'h0008;
		rom[44]   	<= 16'h0008;
		rom[45]   	<= 16'h0008;
		rom[46]   	<= 16'h0008;
		rom[47]   	<= 16'h0;
		rom[48]   	<= 16'h0;
		rom[49]   	<= 16'h0;
		rom[50]   	<= 16'h0;
		rom[51]   	<= 16'h0;
		rom[52]   	<= 16'h0;
		rom[53]   	<= 16'h0008;
		rom[54]   	<= 16'h0;
		rom[55]   	<= 16'h0;
		rom[56]   	<= 16'h0;
		rom[57]   	<= 16'h0;
		rom[58]   	<= 16'h0;
		rom[59]   	<= 16'h0;
		rom[60]   	<= 16'h1010;
		rom[61]   	<= 16'h0005;
		rom[62]   	<= 16'h80c7;
		rom[63]   	<= 16'h0004;
		rom[64]   	<= 16'h0007;
		rom[65]   	<= 16'h0;
		rom[66]   	<= 16'h0003;
		rom[67]   	<= 16'h0003;
		rom[68]   	<= 16'h0203;
		rom[69]   	<= 16'h1010;
		rom[70]   	<= 16'h1010;
		rom[71]   	<= 16'h1010;
		rom[72]   	<= 16'h0010;
		rom[73]   	<= 16'h00a8;
		rom[74]   	<= 16'h0010;
		rom[75]   	<= 16'h0028;
		rom[76]   	<= 16'h0010;
		rom[77]   	<= 16'h2020;
		rom[78]   	<= 16'h1010;
		rom[79]   	<= 16'h0014;
		rom[80]   	<= 16'h8000;
		rom[81]   	<= 16'h0007;
		rom[82]   	<= 16'h8000;
		rom[83]   	<= 16'h0007;
		rom[84]   	<= 16'h0008;
		rom[85]   	<= 16'h0;
		rom[86]   	<= 16'h0020;
		rom[87]   	<= 16'h0004;
		rom[88]   	<= 16'h8000;
		rom[89]   	<= 16'h0007;
		rom[90]   	<= 16'h0004;
		rom[91]   	<= 16'h0001;
		rom[92]   	<= 16'h005a;
		rom[93]   	<= 16'h2d13;
		rom[94]   	<= 16'h41ff;
		rom[95]   	<= 16'h231d;
		rom[96]   	<= 16'h0020;
		rom[97]   	<= 16'h0020;
		rom[98]   	<= 16'h0;
		rom[99]   	<= 16'h0020;
		rom[100]   	<= 16'h0020;
		rom[101]   	<= 16'h0;
		rom[102]   	<= 16'h0;
		rom[103]   	<= 16'h0;
		rom[104]   	<= 16'h0;
		rom[105]   	<= 16'h0;
		rom[106]   	<= 16'h0;
		rom[107]   	<= 16'h0;
		rom[108]   	<= 16'h0;
		rom[109]   	<= 16'h0;
		rom[110]   	<= 16'h0;
		rom[111]   	<= 16'h0;
		rom[112]   	<= 16'h0067;
		rom[113]   	<= 16'ha700;
		rom[114]   	<= 16'ha700;
		rom[115]   	<= 16'h0c00;
		rom[116]   	<= 16'h0600;
		rom[117]   	<= 16'h5617;
		rom[118]   	<= 16'h6b75;
		rom[119]   	<= 16'h6b75;
		rom[120]   	<= 16'ha500;
		rom[121]   	<= 16'hab00;
		rom[122]   	<= 16'ha940;
		rom[123]   	<= 16'ha709;
		rom[124]   	<= 16'ha700;
		rom[125]   	<= 16'hff00;
		rom[126]   	<= 16'ha900;
		rom[127]   	<= 16'ha900;
		rom[128]   	<= 16'h0022;
		rom[129]   	<= 16'h1f04;
		rom[130]   	<= 16'h0;
		rom[131]   	<= 16'h1b06;
		rom[132]   	<= 16'h1d08;
		rom[133]   	<= 16'h0;
		rom[134]   	<= 16'h1806;
		rom[135]   	<= 16'h1a08;
		rom[136]   	<= 16'h0;
		rom[137]   	<= 16'h0;
		rom[138]   	<= 16'h0;
		rom[139]   	<= 16'h0;
		rom[140]   	<= 16'h0;
		rom[141]   	<= 16'h0;
		rom[142]   	<= 16'h0;
		rom[143]   	<= 16'h0;
		rom[144]   	<= 16'h07d0;
		rom[145]   	<= 16'h0;
		rom[146]   	<= 16'h0001;
		rom[147]   	<= 16'h0;
		rom[148]   	<= 16'h0;
		rom[149]   	<= 16'h0;
		rom[150]   	<= 16'h0;
		rom[151]   	<= 16'h0;
		rom[152]   	<= 16'h0;
		rom[153]   	<= 16'h0;
		rom[154]   	<= 16'h0;
		rom[155]   	<= 16'h0;
		rom[156]   	<= 16'h0;
		rom[157]   	<= 16'h0;
		rom[158]   	<= 16'h0;
		rom[159]   	<= 16'h0;
		rom[160]   	<= 16'h0;
		rom[161]   	<= 16'h0;
		rom[162]   	<= 16'h0;
		rom[163]   	<= 16'h0;
		rom[164]   	<= 16'h0;
		rom[165]   	<= 16'h0;
		rom[166]   	<= 16'h0;
		rom[167]   	<= 16'h0;
		rom[168]   	<= 16'h0;
		rom[169]   	<= 16'h0;
		rom[170]   	<= 16'h0;
		rom[171]   	<= 16'h0;
		rom[172]   	<= 16'h0;
		rom[173]   	<= 16'h0;
		rom[174]   	<= 16'h0020;
		rom[175]   	<= 16'h0;
		rom[176]   	<= 16'h0;
		rom[177]   	<= 16'h0;
		rom[178]   	<= 16'h0;
		rom[179]   	<= 16'h0;
		rom[180]   	<= 16'h0;
		rom[181]   	<= 16'h0;
		rom[182]   	<= 16'h0;
		rom[183]   	<= 16'h0;
		rom[184]   	<= 16'h0;
		rom[185]   	<= 16'h0;
		rom[186]   	<= 16'h0;
		rom[187]   	<= 16'h0;
		rom[188]   	<= 16'h0;
		rom[189]   	<= 16'h0;
		rom[190]   	<= 16'h0;
		rom[191]   	<= 16'h0;
		rom[192]   	<= 16'h0;
		rom[193]   	<= 16'h0;
		rom[194]   	<= 16'h0;
		rom[195]   	<= 16'h0;
		rom[196]   	<= 16'h0;
		rom[197]   	<= 16'h0;
		rom[198]   	<= 16'h0;
		rom[199]   	<= 16'h0;
		rom[200]   	<= 16'h0;
		rom[201]   	<= 16'h0;
		rom[202]   	<= 16'h0;
		rom[203]   	<= 16'h0;
		rom[204]   	<= 16'h0;
		rom[205]   	<= 16'h0;
		rom[206]   	<= 16'h0;
		rom[207]   	<= 16'h0;
		rom[208]   	<= 16'h0;
		rom[209]   	<= 16'h0;
		rom[210]   	<= 16'h0;
		rom[211]   	<= 16'h0;
		rom[212]   	<= 16'h0;
		rom[213]   	<= 16'h0;
		rom[214]   	<= 16'h0;
		rom[215]   	<= 16'h0;
		rom[216]   	<= 16'h0;
		rom[217]   	<= 16'h0;
		rom[218]   	<= 16'h0;
		rom[219]   	<= 16'h0;
		rom[220]   	<= 16'h0;
		rom[221]   	<= 16'h0;
		rom[222]   	<= 16'h0;
		rom[223]   	<= 16'h0;
		rom[224]   	<= 16'h0;
		rom[225]   	<= 16'h0;
		rom[226]   	<= 16'h0;
		rom[227]   	<= 16'h0;
		rom[228]   	<= 16'h0;
		rom[229]   	<= 16'h0;
		rom[230]   	<= 16'h0;
		rom[231]   	<= 16'h0;
		rom[232]   	<= 16'h0;
		rom[233]   	<= 16'h0;
		rom[234]   	<= 16'h0;
		rom[235]   	<= 16'h0;
		rom[236]   	<= 16'h0;
		rom[237]   	<= 16'h0;
		rom[238]   	<= 16'h0;
		rom[239]   	<= 16'h0;
		rom[240]   	<= 16'h0;
		rom[241]   	<= 16'h0;
		rom[242]   	<= 16'h0;
		rom[243]   	<= 16'h0;
		rom[244]   	<= 16'h0;
		rom[245]   	<= 16'h0;
		rom[246]   	<= 16'h0;
		rom[247]   	<= 16'h0;
		rom[248]   	<= 16'h0;
		rom[249]   	<= 16'h0;
		rom[250]   	<= 16'h0;
		rom[251]   	<= 16'h0;
		rom[252]   	<= 16'h0;
		rom[253]   	<= 16'h0;
		rom[254]   	<= 16'h0;
		rom[255]   	<= 16'h1801;
end

endmodule
